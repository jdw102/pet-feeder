module and_op(
    input[31:0] A, B,
    output[31:0] out
    );
    and a0(out[0], A[0], B[0]);
    and a1(out[1], A[1], B[1]);
    and a2(out[2], A[2], B[2]);
    and a3(out[3], A[3], B[3]);
    and a4(out[4], A[4], B[4]);
    and a5(out[5], A[5], B[5]);
    and a6(out[6], A[6], B[6]);
    and a7(out[7], A[7], B[7]);
    and a8(out[8], A[8], B[8]);
    and a9(out[9], A[9], B[9]);
    and a10(out[10], A[10], B[10]);
    and a11(out[11], A[11], B[11]);
    and a12(out[12], A[12], B[12]);
    and a13(out[13], A[13], B[13]);
    and a14(out[14], A[14], B[14]);
    and a15(out[15], A[15], B[15]);
    and a16(out[16], A[16], B[16]);
    and a17(out[17], A[17], B[17]);
    and a18(out[18], A[18], B[18]);
    and a19(out[19], A[19], B[19]);
    and a20(out[20], A[20], B[20]);
    and a21(out[21], A[21], B[21]);
    and a22(out[22], A[22], B[22]);
    and a23(out[23], A[23], B[23]);
    and a24(out[24], A[24], B[24]);
    and a25(out[25], A[25], B[25]);
    and a26(out[26], A[26], B[26]);
    and a27(out[27], A[27], B[27]);
    and a28(out[28], A[28], B[28]);
    and a29(out[29], A[29], B[29]);
    and a30(out[30], A[30], B[30]);
    and a31(out[31], A[31], B[31]);
endmodule